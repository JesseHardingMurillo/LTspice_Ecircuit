*FULL wave circuit with Diode
*------------------------------------------------------------------------------------------------------------------------------------------
*Circuit
*------------------------------------------------------------------------------------------------------------------------------------------
V1	IN 		0 		SINE	({p_offset} {p_ampl} {p_freq})
D1 	OUT_N 	IN 		{Dmodel} ; Cambiar out_p y out_n
D2 	IN 		OUT_P 	{Dmodel}
D3 	OUT_N 	0 		{Dmodel}
D4 	0 		OUT_P 	{Dmodel}
R1 	OUT_P 	OUT_N 	{p_r1}
*------------------------------------------------------------------------------------------------------------------------------------------
*Models
*------------------------------------------------------------------------------------------------------------------------------------------
.model 1 ako:1N4148 						; Silicon
.model 2 ako:1N5817							; Schotty
.model 3 ako:1N5373B 						; Zener
*Standard library
.lib C:\Users\jesse\AppData\Local\LTspice\lib\cmp\standard.dio
*------------------------------------------------------------------------------------------------------------------------------------------
*Parameters: User input
*------------------------------------------------------------------------------------------------------------------------------------------
.param		p_r1			1k 				; Resistor Value
.param		p_n_cycles		5				; Number of cycles
.param		p_offset		0				; Offset
.param		p_ampl			10				; Amplitude
.param		p_freq			10k				; Frequency
*------------------------------------------------------------------------------------------------------------------------------------------
*Parameters: Automatic calculation
*------------------------------------------------------------------------------------------------------------------------------------------
.param		p_period		1/p_freq		; Period
.param		p_start_time	4*p_period		; Start, for measurement's purposes
.param		p_stop_time		5*p_period		; Stop, for measurement's purposes
*------------------------------------------------------------------------------------------------------------------------------------------
*Measurements
*------------------------------------------------------------------------------------------------------------------------------------------
.meas		TRAN	Vin_max			MAX		V(in)				From p_start_time to p_stop_time
.meas		TRAN	Vout_max		MAX		V(out,2)			From p_start_time to p_stop_time
.meas		TRAN	Diff_Vin_Vout	PARAM	Vin_max-Vout_max	; Vmax(in) - Vmax(out)
*------------------------------------------------------------------------------------------------------------------------------------------
* ANALYSIS
*------------------------------------------------------------------------------------------------------------------------------------------
.tran {p_period*p_n_cycles}
.step param Dmodel list 1 2 3
.PLOT
.PROBE
.END
