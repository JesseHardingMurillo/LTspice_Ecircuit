*MUX CIRCUIT
*-----------------------------------------------------------------------------
*NOTES
*-----------------------------------------------------------------------------



*-----------------------------------------------------------------------------
*Parameters: User Input
*-----------------------------------------------------------------------------


*=============================================================================
* Calibration
*=============================================================================




*-----------------------------------------------------------------------------
*Libraries, Models and includes
*-----------------------------------------------------------------------------
.lib ./sub_gates.lib



*-----------------------------------------------------------------------------
*CIRCUIT
*-----------------------------------------------------------------------------
;.SUBCKT NAND 1 2 3 4
* TERMINALS A B OUT VCC


;Vselec1	select0	0 	PWL(9.99m 0 10m 5)
;Vselec2	select1	0 	PWL(9.99m 0 10m 5)

Vselec1	ATB_SEL[0]	0	1
Vselec2	ATB_SEL[1]	0 	1

Vin0	in[0]		0	0v
Vin1 	in[1]		0	1V
Vin2	in[2]		0	2v
Vin3 	in[3]		0   3V

.SUBCKT Mux4_1_Behavioral sel[0] sel[1] in[0] in[1] in[2] in[3] OUT
Bmux OUT 0 V={IF(V(sel[0])<1 & V(sel[1])<1, V(in[0]),
+IF(V(sel[0])>=1 & V(sel[1])<1, V(in[1]),
+IF(V(sel[0])<1 & V(sel[1])>=1, V(in[2]),V(in[3]))))}
.ends Mux4_1_Behavioral

XMux4_1 ATB_SEL[0] ATB_SEL[1] in[0] in[1] in[2] in[3] out Mux4_1_Behavioral
*-----------------------------------------------------------------------------
*MEASUREMENTS
*-----------------------------------------------------------------------------


*-----------------------------------------------------------------------------
* SIMULATOR OPTIONS
*-----------------------------------------------------------------------------


*-----------------------------------------------------------------------------
* ANALYSIS
*-----------------------------------------------------------------------------



;.AC 	DEC 	10 	10 	10MEG
.TRAN 	1US  	15m
.PROBE
.END
