ABM_RMS1.CIR
*
V1	1	0	SIN(0V 1V 10KHZ)
R1	1	0	1MEG

*
ESQR	2	0	VALUE = {  V(1)*V(1) }
R2	2	0	1MEG
*
GINT	0	3	VALUE = {  V(2)  }
CINT	3	0	1
R3	3	0	1MEG
*
EAVE	4	0	VALUE = { V(3)/TIME }
R4	4	0	1MEG
*
ESQRT	5	0	VALUE = { SQRT( V(4) ) }
R5	5	0	1MEG
*
*
* ANALYSIS
.TRAN 	1US  200US  UIC
*
* VIEW RESULTS
.PRINT	TRAN 	V(1) V(2) V(4) V(5)
.IC V(1)=0V V(2)=0V V(3)=0V V(4)=0V
.PROBE
.END
