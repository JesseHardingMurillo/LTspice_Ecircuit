ABM_VALUE1.CIR
*
V1	1	0	SIN(0V 1V 10KHZ)
R1	1	0	1K
V2	2	0	SIN(0V 1V 1KHZ)
R2	2	0	1K
V3	3	0	PWL(0US -5V 500US 5V)	; PIECE WISE LINEAR
R3	3	0	1K
*E|G{name} {+node} {-node} VALUE {expression}
ESUM	4	0	VALUE = { (V(1)+V(3))/5 }
R4	4	0	1MEG
EMULT	5	0	VALUE = { 2*V(1)*V(2)}
*EMULT	5	0	VALUE = { 2*V(1)*V(2)*2*v(1) }
R5	5	0	1M
*EGEGEPWR	6	0	VALUE = { ABS(V(1)*	I(V1)) }
EGEGEPWR	6	0	VALUE = { ABS(V(1)* 2 *	I(V1)) }
R6	6	0	1MEG
EDIFF	7	0	VALUE = { TANH(V(3))}
R7	7	0	1MEG
*
* ANALYSIS
.TRAN 	5US  500US
*.Tran 1m
*
* VIEW RESULTS
.PRINT	TRAN 	V(1) V(2) V(3) V(4) V(5) V(6(7)
.PROBE
.END
