OPAMP2.CIR - OPAMP MODEL (LEVEL 2)
*--------------------------------------------------------------------------
*Notes
*--------------------------------------------------------------------------
*                IN+ IN- VCC  VEE OUT
*.SUBCKT OPAMP2   1   2 	 101  102 81

*--------------------------------------------------------------------------
*Circuit
*--------------------------------------------------------------------------
* POWER SUPPLIES
VCC	10	0	DC	5V
VEE	0	11	DC	5V

*Open loop
XOPx1	1 	0  	10 11 out3	OPAMP3
XOPx2	1 	0  	10 11 out4 	OPAMP2
RL	out	0	1K

* SIGNAL SOURCE
VS		1	0	AC 1 SIN(0V  6VPEAK  10KHZ)
;*Inversor
R1i		1	2x		10K
R2i		2x	OUT1	10K
XOP1	0 	2x	10 	11 	OUT1	OPAMP3

*No inversor
R1		2	0		10K
R2		2	OUT2	0.1K
XOP2	1	2	10 	11	OUT2	OPAMP3



*--------------------------------------------------------------------------
*Measurements
*--------------------------------------------------------------------------
.INCLUDE OPAMP_Saturation.meas
*--------------------------------------------------------------------------
*Funtions
*--------------------------------------------------------------------------
.func dB_to_Av(dB)	{10**(db/20)}
.INCLUDE Opmodel2.lib
.INCLUDE Opmodel2_Voltage_limiter.lib


*-----------------------------------------------------------------------------
* SIMULATOR OPTIONS
*-----------------------------------------------------------------------------
;.option meascplxfmt=bode			; default
*.option meascplxfmt=polar
;.option meascplxfmt=cartesian

*--------------------------------------------------------------------------
* ANALYSIS
*--------------------------------------------------------------------------
;.TRAN 	0.1US  5US
;.TRAN 	1m
.AC 	DEC 	10 0.1HZ 10MEGHZ
*
* VIEW RESULTS
;.PRINT	TRAN 	V(out)
;.PRINT	AC 	V(out)
.PROBE
.END
