*NOTE:
*VTH

*Half wave circuit with Diode
*------------------------------------------------------------------------------------------------------------------------------------------
*Circuit
*------------------------------------------------------------------------------------------------------------------------------------------
*Source
VS in	0	AC 1 SIN({p_offset} {p_ampl} {p_freq})
D1 in	0	1N4148
*D1 in	0	1N914
*R1	out	0	{p_r1}
*------------------------------------------------------------------------------------------------------------------------------------------
*Models
*------------------------------------------------------------------------------------------------------------------------------------------
*.model MyIdealDiode  D(1N4148) ;MyIdealDiodeJesse
.model D D
*------------------------------------------------------------------------------------------------------------------------------------------
*Standard library
*------------------------------------------------------------------------------------------------------------------------------------------
.lib C:\Users\jesse\AppData\Local\LTspice\lib\cmp\standard.dio
*------------------------------------------------------------------------------------------------------------------------------------------
*Parameters:User input
*------------------------------------------------------------------------------------------------------------------------------------------
.param p_r1	1k
.param p_offset	0
.param p_ampl	1
.param p_freq	1k
*------------------------------------------------------------------------------------------------------------------------------------------
*Parameters:Measure
*------------------------------------------------------------------------------------------------------------------------------------------
*.MEAS DC Ith Find I(D1) WHEN V(IN)=700mV
.meas DC Vth FIND V(in) WHEN I(D1)=0.0111974
*------------------------------------------------------------------------------------------------------------------------------------------
* ANALYSIS
*------------------------------------------------------------------------------------------------------------------------------------------
.dc Vs 0 2
.step temp -40  180 40
*.tran 30us
.END
