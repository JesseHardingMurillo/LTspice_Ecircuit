OPAMP2.CIR - OPAMP MODEL (LEVEL 2)
*--------------------------------------------------------------------------
*Circuit
*--------------------------------------------------------------------------
* SIGNAL SOURCE
VS	1	0	AC 1	PWL(0US 0V   0.01US 1v  100US 1V)

*
* POWER SUPPLIES
VCC	10	0	DC	+5V
VEE	11	0	DC	-5V

*OP AMP TEST DRIVE
R1	0	2	1 		;	 Open loop

R2	2	out	1		; 	 Feedback (Closed Loop)

XOP	1 	2  10 11 out OPAMP2
*RL	out	0	100K

*--------------------------------------------------------------------------
*Measurements
*--------------------------------------------------------------------------
.INCLUDE OPAMP_INTERMEDIATE.meas
*--------------------------------------------------------------------------
*Funtions
*--------------------------------------------------------------------------
.func dB_to_Av(dB)	{10**(db/20)}
.INCLUDE Opmodel2.lib


*-----------------------------------------------------------------------------
* SIMULATOR OPTIONS
*-----------------------------------------------------------------------------
;.option meascplxfmt=bode			; default
*.option meascplxfmt=polar
;.option meascplxfmt=cartesian

*--------------------------------------------------------------------------
* ANALYSIS
*--------------------------------------------------------------------------
;.TRAN 	0.1US  5US
.TRAN 	0.1US  100US
*.AC 	DEC 	5 0.1HZ 10MEGHZ
*
* VIEW RESULTS
.PRINT	TRAN 	V(out)
.PRINT	AC 	V(out)
.PROBE
.END
