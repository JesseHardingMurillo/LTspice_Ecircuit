SAMPLING.CIR - SAMPLING CIRCUIT
*
VS	1	0	SIN(0VOFF	5VPEAK	1KHZ)
R1	1	0	1MEG
*
* FILTER BLOCK
* NO FILTER
EBUFFER	2 0	1 0	1
R3	2	0	1MEG
*
* 2ND ORDER LP FILTER
*E_LPFILTER 2 0 LAPLACE { V(1) }  {1 / ( (s*s)/(6.28*6.28*10000*10000) + s/(0.707*6.28*10000) + 1) }
*
*
* SAMPLE & HOLD CIRCUIT
S1	2 5	10 0 	SRES	
CH	5	0	0.01UF
RH	5	0	10MEG
*
* S/H CONTROL VOLTAGE
VC1	10	0	PULSE(0V 5V 0US 0.1US 0.1US 1US 50US)
R10	10	0	1MEG
*
*
.MODEL	SRES	VSWITCH(VON=5V VOFF=0V RON=10 ROFF=10MEG)
* 
* ANALYSIS
.TRAN 	1US  	1000US  0US 2US
*
* VIEW RESULTS
.PLOT	TRAN	V(2) V(5)
.PROBE
.END
