*DAC OF 8 BITS
*----------------------------------------------------------------------------
*PARAMETERS
*----------------------------------------------------------------------------
.PARAM Voff				0
.PARAM Vcc				5
.PARAM td				0
.PARAM tt				1n
.PARAM T				1m
.PARAM N_BITS			4
.PARAM quant_step_size 	{((2**N_BITS)-1)/(2**N_BITS )}


*----------------------------------------------------------------------------
*CIRCUIT
*----------------------------------------------------------------------------
*SOURCES
V0 in[0] 0 PULSE({Voff} {Vcc} {T/2} {tt} {tt} {T*1/2} {T*1})
V1 in[1] 0 PULSE({Voff} {Vcc} {T/2*2} {tt} {tt} {T*2/2} {T*2})
V2 in[2] 0 PULSE({Voff} {Vcc} {T/2*4} {tt} {tt} {T*4/2} {T*4})
V3 in[3] 0 PULSE({Voff} {Vcc} {T/2*8} {tt} {tt} {T*8/2} {T*8})

*DAAC
Edac2 out_dac 0 VALUE = { (  (V(in[0])/{Vcc})*1 + (V(in[1])/{Vcc})*2 + (V(in[2])/{Vcc})*4 + (V(in[3])/{Vcc})*8  ) * quant_step_size}

*----------------------------------------------------------------------------
*ANALYSIS
*----------------------------------------------------------------------------
.TRAN 0 8m 0 {15/16/100}
