ADC2bits
*-----------------------------------------------------------------------------
*NOTES
*-----------------------------------------------------------------------------



*-----------------------------------------------------------------------------
*Parameters: User Input
*-----------------------------------------------------------------------------
.param Voff=0
.param Vcc=5
.param td=0
.param tt=1n
.param T=1m
*=============================================================================
* Calibration
*=============================================================================


*-----------------------------------------------------------------------------
*Libraries, Models and includes
*-----------------------------------------------------------------------------
.LIB SAMPLE_HOLD.lib


*-----------------------------------------------------------------------------
*CIRCUIT
*-----------------------------------------------------------------------------
Vs	in 	0	PWL file=Wave_Input.txt
Vclk clk 0 PULSE( {Voff} {Vcc}  {T/4} {tt} {tt} {T*1/2/2} {T*1/2})

;.SUBCKT SAMPLE_HOLD IN 	CLK OUT
Xsample in clk out SAMPLE_HOLD


*-----------------------------------------------------------------------------
*MEASUREMENTS
*-----------------------------------------------------------------------------


*-----------------------------------------------------------------------------
* SIMULATOR OPTIONS
*-----------------------------------------------------------------------------


*-----------------------------------------------------------------------------
* ANALYSIS
*-----------------------------------------------------------------------------



;.AC 	DEC 	10 	10 	10MEG
.TRAN 	1US  	3m
.PROBE
.END
