LOGIC_SW.CIR - BASIC LOGIC GATES USING SWITCHES
*----------------------------------------------------------------------------
*Observations
*----------------------------------------------------------------------------
*La NAND se apaga cuando cuando VA Y VB se hace 1
*La NOR presenta un peque�o pico cuando se  VA esta bajando y vB subiendo
*Los mismo que para en la NOR, pasa en la Or

*----------------------------------------------------------------------------
*Circuit
*----------------------------------------------------------------------------
VCC	10	0	5V
* INPUT A AND B, COUNT IN BINARY 0 - 3
*			PULSE( {v1} {v2} {tdelay} {trise} {tfall} {width} {period} )
VA	1	0	PULSE(5V 0V 0NS 10NS 10NS 90NS 200NS)
VB	2	0	PULSE(5V 0V 0NS 10NS 10NS 190NS 400NS)
VC	11	0	PULSE(5V 0V 0NS 10NS 10NS 290NS 800NS)

*----------------------------------------------------------------------------
*Gates
XNAND1	1 2 3 	10	NAND	; 2 inputs
*XNOR1 	1 2 3 	10 	NOR
*XNOT1 	1 3 10 		NOT
*XAND1 	1 2 3 	10 	AND
*XOR1 	1 2 3 	10 	OR
*XNAND2  1 2 11	3	10 	NAND3	; 3 inputs
*xor	1 2 3	10	XOR
*----------------------------------------------------------------------------
* LOGIC GATE SUBCIRCUITS
*----------------------------------------------------------------------------
.include sub_gates.lib

*----------------------------------------------------------------------------
* ANALYSIS
*----------------------------------------------------------------------------
.TRAN 	5NS  	400NS
*
* VIEW RESULTS
.PRINT	TRAN 	V(1) V(2) V(11) V(3)
.PROBE
.END
