*Half wave circuit with Diode
*------------------------------------------------------------------------------------------------------------------------------------------
*Circuit
*------------------------------------------------------------------------------------------------------------------------------------------
*Source
VS in	0	AC 1 SIN({p_offset} {p_ampl} {p_freq})
*D1 in	out	1N5817	;Vd ~ 100mV , Vreverse ~ -32.4 mV
D1 in	out	1N4148
R1	out	0	{p_r1}
*------------------------------------------------------------------------------------------------------------------------------------------
*Models
*------------------------------------------------------------------------------------------------------------------------------------------
*.model MyIdealDiode  D(1N4148) ;MyIdealDiodeJesse
.model D D
*------------------------------------------------------------------------------------------------------------------------------------------
*Standard library
*------------------------------------------------------------------------------------------------------------------------------------------
.lib C:\Users\jesse\AppData\Local\LTspice\lib\cmp\standard.dio
*------------------------------------------------------------------------------------------------------------------------------------------
*Parameters:User input
*------------------------------------------------------------------------------------------------------------------------------------------
.param p_r1	1k
.param p_offset	0
.param p_ampl	1
.param p_freq	1k
*------------------------------------------------------------------------------------------------------------------------------------------
* ANALYSIS
*------------------------------------------------------------------------------------------------------------------------------------------
*.AC 	DEC 	5 1 500MEG
.tran 10ms
.PLOT
.PROBE
.END
