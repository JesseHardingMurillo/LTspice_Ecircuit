ADC2bits
*-----------------------------------------------------------------------------
*NOTES
*-----------------------------------------------------------------------------



*-----------------------------------------------------------------------------
*Parameters: User Input
*-----------------------------------------------------------------------------
.param vhigh 1
.param vlow 0
.param vref 15

*=============================================================================
* Calibration
*=============================================================================




*-----------------------------------------------------------------------------
*Libraries, Models and includes
*-----------------------------------------------------------------------------
* Subcircuito para un ADC de 2 bits
.subckt ADC_2bit in out[1] out[0] vdac[1] vdac[0]
B1_vdac vdac[1] 0 V=vref * (Vhigh/2 + Vlow/4)
*B1_out  out[1]  0 V= V(in)>=V(vdac[1]) ? vhigh : vlow
B1_out  out[1]  0 V= {V(in)/((2**2) - 1)}>=V(vdac[1]) ? vhigh : vlow

B0_vdac vdac[0] 0 V=vref * (V(out[1])/2 + Vhigh/4)
*B0_out  out[0]  0 V= V(in)>=V(vdac[0]) ? vhigh : vlow
B0_out  out[0]  0 V= {V(in)/((2**2) - 1)}>=V(vdac[0]) ? vhigh : vlow

*Carry OUT8

.ends

*-----------------------------------------------------------------------------
* Subcircuito para un ADC de 4bits
.subckt ADC_4bit in out[3] out[2] out[1] out[0]
B3_vdac vdac[3] 0 V= vref * (vhigh/2 + vlow/4 + vlow/8 + vlow/16)
B3_out  out[3]  0 V= V(in)>=V(vdac[3]) ? vhigh : vlow


B2_vdac vdac[2] 0 V=vref * (V(out[3])/2 + vhigh/4 + vlow/8 + vlow/16)
B2_out  out[2]  0 V= V(in)>=V(vdac[2]) ? vhigh : vlow

B1_vdac vdac[1] 0 V=vref * (V(out[3])/2 + V(out[2])/4 + vhigh/8 + vlow/16)
B1_out  out[1]  0 V= V(in)>=V(vdac[1]) ? vhigh : vlow


B0_vdac vdac[0] 0 V=vref * (V(out[3])/2 + V(out[2])/4 + V(out[1])/8 + vhigh/16)
B0_out  out[0]  0 V= V(in)>=V(vdac[0]) ? vhigh : vlow
.ends

*-----------------------------------------------------------------------------
*CIRCUIT
*-----------------------------------------------------------------------------
V1 in 0 11

;XDac_4bits in out1[3] out1[2] out1[1] out1[0] ADC_4bit

XDac_2bits1 in out1[1] out1[0] dac1[1] dac1[0] ADC_2bit

;XDac_2bits2 in out2[1] out3[0] ADC_2bit
*-----------------------------------------------------------------------------
*MEASUREMENTS
*-----------------------------------------------------------------------------


*-----------------------------------------------------------------------------
* SIMULATOR OPTIONS
*-----------------------------------------------------------------------------


*-----------------------------------------------------------------------------
* ANALYSIS
*-----------------------------------------------------------------------------



;.AC 	DEC 	10 	10 	10MEG
.TRAN 	1US  	1m
.PROBE
.END
