OP_BANDWIDTH1.CIR - OPAMP BANDWIDTH
*
VS	1	0	AC 1V	PWL(0US 0V   0.01US 1V  100US 1V)
*
*
* NON-INVERTING AMPLIFIER
R1	2	0	10K
R2	2	4	10K
XOP1	1 2	4	OPAMP1
*
* INVERTING AMPLIFIER
R_1	1	12	10K
R_2	12	14	10K
XOP2	0 12	14	OPAMP1
*
*
* OPAMP MACRO MODEL, SINGLE-POLE
* connections:      non-inverting input
*                   |   inverting input
*                   |   |   output
*                   |   |   |
.SUBCKT OPAMP1      1   2   6
* INPUT IMPEDANCE
RIN	1	2	10MEG
* DCGAIN =100K AND POLE1=1/(2*PI*RP1*CP1)=100HZ
* GBP = DCGAIN X POLE1 = 10MHZ
EGAIN	3 0	1 2	100K
RP1	3	4	1000
CP1	4	0	1.5915UF
* OUTPUT BUFFER AND RESISTANCE
EBUFFER	5 0	4 0	1
ROUT	5	6	10
.ENDS
*
*
* ANALYSIS
.AC 	DEC 	5 10 100MEG
*.TRAN 	0.01US  0.5US
*
* VIEW RESULTS
*.PRINT	AC 	VM(4)
*.PRINT	TRAN 	V(4) V(14)
.PROBE
.END
