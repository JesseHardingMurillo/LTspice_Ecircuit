HighPassFilter
*-----------------------------------------------------------------------------
*NOTES
*-----------------------------------------------------------------------------
* This a LPF for replace with a step

*-----------------------------------------------------------------------------
*Libraries, Models and includes
*-----------------------------------------------------------------------------
.LIB HPF.LIB

*=============================================================================
* Calibration
*=============================================================================
.PARAM C 	5n
.PARAM fc 	5k


*-----------------------------------------------------------------------------
*CIRCUIT
*-----------------------------------------------------------------------------
*
VS	1	0	AC 1 SIN(0VOFF 1VPEAK 2KHZ)
*
XHPF 1 OUT HPF	PARAMS: C = {C}	fc = {fc}

*-----------------------------------------------------------------------------
* ANALYSIS
*-----------------------------------------------------------------------------
.AC 	DEC 	10 	10 	10MEG
.PROBE
.END
