OPFIL1.CIR - RC LOW-PASS FILTER WITH OPAMP BUFFER
*----------------------------------------------------------------------------
*NOTES
*----------------------------------------------------------------------------




*-----------------------------------------------------------------------------
*FUNTIONS
*-----------------------------------------------------------------------------
.func cal_Xc(Freq,C) 	{-1/(2*pi*Freq*C)}
.func Vec_Mag(A,B)		{sqrt(A**2+B**2)}
.func Vec_angle(A,B)	{atan(A/B)}
.func AvtodB(Av)		{20*(log10(Av))}
.func dBtoAv(dB)		{10**(dB/20)}


*----------------------------------------------------------------------------
*PARAMETERS: USER INPUT
*----------------------------------------------------------------------------
.PARAM p_Vs 1

.PARAM p_R1 15.9K
.PARAM p_C1	1000pF

.PARAM p_Ra 100MEG
.PARAM p_Rb 1k

*----------------------------------------------------------------------------
*PARAMETERS: AUTOMATIC CALCULATION
*----------------------------------------------------------------------------

*----------------------------------------------------------------------------
*Circuit
*----------------------------------------------------------------------------
* SINGLE POLE
*
VS	IN	0	AC	{p_Vs}
*
R1	IN	2		{p_R1}
C1	2	0		{p_C1}
*
* UNITY GAIN AMPLIFIER, RA=OPEN, RB=SHORT
RA	4	0		{p_Ra}
RB	4	OUT		{p_Rb}
XOP	2 	4	OUT	OPAMP1

*----------------------------------------------------------------------------
*Mesurments
*---------------------------------------------------------------------------
.INCLUDE LPF_OPAMP.MEAS

*----------------------------------------------------------------------------
*Subcircuit
*---------------------------------------------------------------------------
* OPAMP MACRO MODEL, SINGLE-POLE
* connections:      non-inverting input
*                   |   inverting input
*                   |   |   output
*                   |   |   |
.SUBCKT OPAMP1	     1   2   6
* INPUT IMPEDANCE
RIN	1	2	10MEG
* DC GAIN (100K) AND POLE 1 (100HZ)
* GBWP = 10MHz
EGAIN   3 0     1 2     100K
RP1     3       4       1K
CP1     4       0       1.5915UF
* OUTPUT BUFFER AND RESISTANCE
EBUFFER 5 0     4 0     1
ROUT    5       6       10
.ENDS
*


*-----------------------------------------------------------------------------
* SIMULATOR OPTIONS
*-----------------------------------------------------------------------------
*.option meascplxfmt=bode			; default
*.option meascplxfmt=polar
.option meascplxfmt=cartesian

*-----------------------------------------------------------------------------
* ANALYSIS
*-----------------------------------------------------------------------------
.AC 	DEC 	10 100 1MEG
.PROBE
.END
