adc_converter
*-----------------------------------------------------------------------------
*NOTES
*-----------------------------------------------------------------------------


*-----------------------------------------------------------------------------
*Parameters: User Input
*-----------------------------------------------------------------------------
.PARAM p_Vdd 15
.PARAM vthreshold 1
.PARAM N_BITS 			8			; Number of bits | FIXED VALUE
.PARAM N_QUANT_LEVELS 	{2**N_BITS}	; Number of Discrete Quantization Levels
.PARAM QUANT_STEP 		{p_Vdd/N_QUANT_LEVELS}
*=============================================================================
* Calibration
*=============================================================================



*-----------------------------------------------------------------------------
*Libraries, Models and includes
*-----------------------------------------------------------------------------
.LIB ADC_SAR.LIB
.LIB DAC.LIB


*-----------------------------------------------------------------------------
*CIRCUIT
*-----------------------------------------------------------------------------
;SOURCES
Vin in 	0 PWL(0 0 20 20)
;Vin in 	0 14.99
Vdd VDD 0 {p_Vdd}				; Fullscale

*/////////////////////////////////////////////////////////////////////////////
;8 BITS ADC SUBCIRCUIT
XADC_SAR_8bits_1 in vdd 0  out[23] out[22] out[21] out[20] out[19] out[18] out[17] out[16] ADC_SAR_8bits_V2 ;MSB

*-----------------------------------------------------------------------------
Xscaler8bits_1 in VDD in_ADC2	 ADCscaler
+N_QUANT_LEVELS	=	{N_QUANT_LEVELS}
+QUANT_STEP 	= 	{QUANT_STEP}

XADC_SAR_8bitsV2 in_ADC2 vdd 0  out[15] out[14] out[13] out[12] out[11] out[10] out[9] out[8] ADC_SAR_8bits_V2

*-----------------------------------------------------------------------------
Xscaler8bits_2 in_ADC2 VDD in_ADC3	 ADCscaler
+N_QUANT_LEVELS	=	{N_QUANT_LEVELS}
+QUANT_STEP 	= 	{QUANT_STEP}

XADC_SAR_8bitsV3 in_ADC3 vdd 0  out[7] 	out[6] out[5] 	out[4] out[3] 	out[2] out[1] out[0] ADC_SAR_8bits_V2 ; LSB
*-----------------------------------------------------------------------------



*-----------------------------------------------------------------------------
*MEASUREMENTS
*-----------------------------------------------------------------------------
;.INCLUDE ADC_SAR_MEASURMENTS.meas


*-----------------------------------------------------------------------------
* SIMULATOR OPTIONS
*-----------------------------------------------------------------------------


*-----------------------------------------------------------------------------
* ANALYSIS
*-----------------------------------------------------------------------------
.TRAN 0 16 0 {15/256/10}
.PROBE
.END
