OP_LIMITER0.CIR - BASIC DIODE LIMITER
*
VS	1	0	SIN(0VDC 10VPEAK 1KHZ)
*
* INVERTING AMPLIFIER
R1	1	2	10K
R2	2	3	1000K
* DIODE LIMITING
*D1	2	3	D1N759
D1	2	3	D1N746
D2	4	3	D1N746

* OP AMP
XOP1	0 2	3	OPAMP1
*
* ZENER DIODES
.model D1N746 D(Is=5u Rs=14 Bv=2.81 Ibv=5u)
.model D1N752 D(Is=0.5u Rs=6 Bv=5.20 Ibv=0.5u)
.model D1N758 D(Is=0.05u Rs=9 Bv=9.49 Ibv=0.05u)
.model D1N759 D(Is=0.05u Rs=12 Bv=12.1 Ibv=0.05u)
*
*
* OPAMP MACRO MODEL, SINGLE-POLE
* connections:      non-inverting input
*                   |   inverting input
*                   |   |   output
*                   |   |   |
.SUBCKT OPAMP1      1   2   6
* INPUT IMPEDANCE
RIN	1	2	10MEG
* DCGAIN =100K AND POLE1=100HZ
* GBP = DCGAIN X POLE1 = 10MHZ
EGAIN	3 0	1 2	100K
RP1	3	4	1000
CP1	4	0	1.5915UF
* OUTPUT BUFFER AND RESISTANCE
EBUFFER	5 0	4 0	1
ROUT	5	6	10
.ENDS
*
*
* ANALYSIS
.TRAN 	10US  2000US
.PROBE
.END
