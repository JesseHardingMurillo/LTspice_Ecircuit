OPFIL1.CIR - RC LOW-PASS FILTER WITH OPAMP BUFFER 
* SINGLE POLE
*
VS	1	0	AC	1
*
R1	1	2	15.9K
C1	2	0	1000PF
*
* UNITY GAIN AMPLIFIER, RA=OPEN, RB=SHORT
RA	4	0	100MEG
RB	4	5	1k
XOP	2 4	5	OPAMP1
*
* OPAMP MACRO MODEL, SINGLE-POLE 
* connections:      non-inverting input
*                   |   inverting input
*                   |   |   output
*                   |   |   |
.SUBCKT OPAMP1	     1   2   6
* INPUT IMPEDANCE
RIN	1	2	10MEG
* DC GAIN (100K) AND POLE 1 (100HZ)
* GBWP = 10MHz
EGAIN   3 0     1 2     100K
RP1     3       4       1K
CP1     4       0       1.5915UF
* OUTPUT BUFFER AND RESISTANCE
EBUFFER 5 0     4 0     1
ROUT    5       6       10
.ENDS
* 
* ANALYSIS
.AC 	DEC 	10 100 1MEG
.PROBE
.END