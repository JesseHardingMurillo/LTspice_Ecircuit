ABM_LAPLACE1.CIR
*
* AC AND STEP INPUT
VS	1	0	AC	1V 	PWL(0US 0V   1US 1V   100US 1V)
R1	1	0	1MEG
*
E_LP_1ST 2 0 LAPLACE { V(1) }  {1 / (s/6280 + 1)}
R2	2	0	1MEG
*E_LP_2ND 3 0 LAPLACE { V(1) }  {1 / ( (s*s)/(6280*6280) + s/(0.707*6280) + 1) }
E_LP_2ND 3 0 LAPLACE { V(1) }  {1 / ( (s*s)/(6280*6280) + s/(0.707*6280) + 1) }
R3	3	0	1MEG
*
* ANALYSIS
*.TRAN 	0.05MS  2.5MS
.AC	DEC 10 100	100K
*
* VIEW RESULTS
.PRINT	TRAN 	V(1) V(2) V(3)
.PRINT	AC	V(2) V(3)
.PROBE
.END
