OPINT.CIR - OPAMP INTEGRATOR
*
* CONTROL VOLTAGE FOR S1
VRESET	4	0	PULSE(0V 5V 0 0.1US 0.1US 100US 110US)
R4	4	0	1MEG
*
* INPUT VOLTAGE
VS	1	0	DC	-1
*
R1	1	2	10K
C1	2	3	1000PF
S1	2 3	4 0 	SRES
XOP	0 2	3	OPAMP1
*
.MODEL	SRES	VSWITCH(VON=0 VOFF=5 RON=100 ROFF=10MEG)
*
* OPAMP MACRO MODEL, SINGLE-POLE
* connections:      non-inverting input
*                   |   inverting input
*                   |   |   output
*                   |   |   |
.SUBCKT OPAMP1      1   2   6
* INPUT IMPEDANCE
RIN	1	2	10MEG
* GAIN BW PRODUCT = 10MHZ = DCGAIN x POLE1
* DC GAIN (100K) AND POLE 1 (100HZ)
EGAIN	3 0	1 2	100K
RP1	3	4	1K
CP1	4	0	1.5915UF
* OUTPUT BUFFER AND RESISTANCE
EOUT	5 0	4 0	1
ROUT	5	6	10
.ENDS
*
* ANALYSIS
.TRAN 	1US  	220US
* VIEW RESULTS
.PLOT	TRAN	V(1) V(3)
*.PRINT	TRAN V(1) V(3)
.PROBE
.END
