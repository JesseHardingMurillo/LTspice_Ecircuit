LPFILTER.CIR - SIMPLE RC LOW-PASS FILTER
*------------------------------------------------------------------------------------------------------------------------------------------
*Circuit
*------------------------------------------------------------------------------------------------------------------------------------------
VS	in	0		AC			1		SIN({p_offset}	{p_amplt}	{p_f})
R1	in	out		{p_r1}
C1	out	0		{p_c1}
*------------------------------------------------------------------------------------------------------------------------------------------
*Parameters
*------------------------------------------------------------------------------------------------------------------------------------------
.param		p_offset		0
.param		p_amplt			1
.param		p_f 			2k
.param		p_r1 			1k
.param		p_c1			0.032UF

.param		p_c_end 		100Khz
*------------------------------------------------------------------------------------------------------------------------------------------
*Measures
.meas 	AC 	Vout_avg		AVG 	V(out)
.meas 	AC 	Vout_max		MAX 	V(out)	FROM p_c_start To p_c_end
.meas	AC 	Vout_min		MIN 	V(out)	FROM p_c_start To p_c_end
.meas 	AC 	Vout_Hz FIND 	V(out) 	at 5khz
*------------------------------------------------------------------------------------------------------------------------------------------
* ANALYSIS
*------------------------------------------------------------------------------------------------------------------------------------------
*DEC, OCT indicate the number of step octal 8 to 8, DEC 10 TO 10
*Complex number format of .meas statement results. One of "polar", "cartesian", or "bode".
.opt	meascplxfmt= cartesian
*ac <oct, dec, lin> <Nsteps> <StartFreq> <EndFreq>
.AC		oct		4		8		10MEG
.PROBE
.END
