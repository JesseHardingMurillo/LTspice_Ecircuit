Inverter Circuit With Gain=2
*----------------------------------------------------------------------------------------------------
*Circuit
*----------------------------------------------------------------------------------------------------
V_VIN	IN	0	AC	1 SIN({p_Voff} {p_Vpeak} {p_Vfreq})		; Vin

Rin		2   IN 		{p_Rref}

X_LM741	0 	2 	VCC	VEE OUT LM741 			; LM741 CL

V_V1    0 	VEE 	{P_V1}
V_V2    VCC 0 		{P_V2}


RRef   	2   OUT		{cal_Rin}
RL		OUT	0		{p_Rl}

*----------------------------------------------------------------------------------------------------
*Parameters: User input
*----------------------------------------------------------------------------------------------------
.PARAM p_Voff 	0
.PARAM p_Vpeak 	5
.PARAM p_Vfreq 	1khz

.PARAM P_V1		5
.PARAM P_V2		5

*PORQUE SE LA CARGA BAJA DE VUELVE CUADRADA
.PARAM p_Rl		1k


.PARAM Gain		1
.PARAM p_Rref	10k

.PARAM p_n_period 3


*----------------------------------------------------------------------------------------------------
*Parameters: Automatic Calculation
*----------------------------------------------------------------------------------------------------
.PARAM cal_Rin 	{Gain*p_Rref}
.PARAM p_period {p_n_period * 1/p_Vfreq}

*----------------------------------------------------------------------------------------------------
*LIBRARIES
*----------------------------------------------------------------------------------------------------
.LIB C:\Users\jesse\OneDrive - Universidad T�cnica Nacional\Cursos Actuales\Proyecto Electronico\MODELS\LM741\lm741.lib

*----------------------------------------------------------------------------------------------------
*Measurements
*----------------------------------------------------------------------------------------------------
.INCLUDE LM741.MEAS

*----------------------------------------------------------------------------------------------------
*Analysis directives
*----------------------------------------------------------------------------------------------------
.TRAN  0 {p_period}
