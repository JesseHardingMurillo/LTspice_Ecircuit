adc_converter
*-----------------------------------------------------------------------------
*NOTES
*-----------------------------------------------------------------------------


*-----------------------------------------------------------------------------
*Parameters: User Input
*-----------------------------------------------------------------------------
.PARAM p_Vdd 15
.PARAM vthreshold 1
.PARAM N_BITS 			4			; Number of bits | FIXED VALUE
.PARAM N_QUANT_LEVELS 	{2**N_BITS}	; Number of Discrete Quantization Levels
.PARAM QUANT_STEP 		{p_Vdd/N_QUANT_LEVELS}
*=============================================================================
* Calibration
*=============================================================================



*-----------------------------------------------------------------------------
*Libraries, Models and includes
*-----------------------------------------------------------------------------
.LIB ADC_SAR.LIB
.LIB DAC.LIB


*-----------------------------------------------------------------------------
*CIRCUIT
*-----------------------------------------------------------------------------
;SOURCES
Vin in 	0 PWL(0 0 20 20)
;Vin in 	0 14.99
Vdd VDD 0 {p_Vdd}				; Fullscale

*/////////////////////////////////////////////////////////////////////////////

;8 BITS INDIVIDUAL PARTS
;XADC_MSB in vdd 0 out[7] out[6] out[5] out[4] ADC_SAR_4bits  ; Working
*-----------------------------------------------------------------------------
;Xscaler8bits in  in_LSB	 ADCscaler
;+N_QUANT_LEVELS	=	{N_QUANT_LEVELS}
;+QUANT_STEP 	= 	{QUANT_STEP}
*-----------------------------------------------------------------------------
;XADC_LSB in_LSB vdd 0 out[3] out[2] out[1] out[0] ADC_SAR_4bits

*/////////////////////////////////////////////////////////////////////////////

;8 BITS ADC SUBCIRCUIT
;XADC_SAR_8bits in vdd vss  out[7] out[6] out[5] out[4] out[3] out[2] out[1] out[0] ADC_SAR_8bits
*-----------------------------------------------------------------------------
; 8 BITS DAC
;E_dac	DAC_OUT	0  value={((1*V(out[0]))+2*V(out[1])+4*V(out[2])+8*V(out[3])+16*V(out[4])+32*V(out[5])+64*V(out[6])+128*V(out[7]))*(V(VDD)/2**(N_BITS*2))}

*/////////////////////////////////////////////////////////////////////////////

;8 BITS ADC SUBCIRCUIT
XADC_SAR_8bitsV2 in vdd 0  out[7] out[6] out[5] out[4] out[3] out[2] out[1] out[0] ADC_SAR_8bits_V2
*-----------------------------------------------------------------------------
; 8 BITS DAC SUBBCIRCUIT
XDAC out[7] out[6] out[5] out[4] out[3] out[2] out[1] out[0] VDD OUT_DAC DAC_8bits


*-----------------------------------------------------------------------------
*MEASUREMENTS
*-----------------------------------------------------------------------------
.INCLUDE ADC_SAR_MEASURMENTS.meas


*-----------------------------------------------------------------------------
* SIMULATOR OPTIONS
*-----------------------------------------------------------------------------


*-----------------------------------------------------------------------------
* ANALYSIS
*-----------------------------------------------------------------------------
.TRAN 0 16 0 {15/256/10}
.PROBE
.END
