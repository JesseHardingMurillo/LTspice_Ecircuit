OPDFR.CIR - OPAMP DIFFERENTIATOR
*
* TRAPEZOIDAL WAVE
VS1	1	0	PULSE(0V 1V 0 10MS 10MS 10MS 40MS)
* SINEWAVE
*VS2	1	0	SIN(0VOFF 1VPEAK 20HZ)
* 1 VRMS FOR AC ANALYSIS
*VS3	1	0	AC	1
*
C1	1	2	10NF
R1	2	3	5K
R2	3	4	500K
XOP	0 3	4	OPAMP1
*
*
* OPAMP MACRO MODEL, SINGLE-POLE
* connections:      non-inverting input
*                   |   inverting input
*                   |   |   output
*                   |   |   |
.SUBCKT OPAMP1      1   2   6
* INPUT IMPEDANCE
RIN	1	2	10MEG
* DCGAIN =100K AND POLE1=1/(2*PI*RP1*CP1)=100HZ
* GBP = DCGAIN X POLE1 = 10MHZ
EGAIN	3 0	1 2	100K
RP1	3	4	1000
CP1	4	0	1.5915UF
* OUTPUT BUFFER AND RESISTANCE
EBUFFER	5 0	4 0	1
ROUT	5	6	10
.ENDS
*
* ANALYSIS
.TRAN 	1MS  100MS
*
* VIEW RESULTS
.PROBE
.END
