ABM_FREQ1.CIR
*
V1	1	0	AC	1V 	PWL(0US 0V  1US 1V  100US 1V  101US 0V  200US 0V )
R1	1	0	1MEG
*
E_LP_FIL 2 0 FREQ {V(1)} (1KHZ, 0DB, 0DEG) (10KHZ, -3DB, -45DEG)  (1000KHZ, -20DB, -90DEG)
R2	2	0	1MEG
E_HP_FIL 3 0 FREQ {V(1)} (1HZ, -40DB, +90DEG) (10KHZ, -3DB, +45DEG)  (100KHZ, 0DB, 0DEG)
R3	3	0	1MEG
*
* ANALYSIS
;.TRAN 	1US  200US
.AC	DEC 5 100	1000K
*
* VIEW RESULTS
.PRINT	TRAN 	V(2) V(3)
.PRINT	AC	V(2) V(3)
.PROBE
.END
