adc_converter
*-----------------------------------------------------------------------------
*NOTES
*-----------------------------------------------------------------------------
* ADC de 24 bits en LTspice con Bus de Salida (0-23) y Full Scale de 15V


*-----------------------------------------------------------------------------
*Parameters: User Input
*-----------------------------------------------------------------------------
.param p_Vfullscale 	15
.param p_resolution 	2		; Number of bits
.param slope			{p_Vfullscale/((2**p_resolution)-1)}


.param FS = 15  ; Full Scale, puedes cambiar este valor seg�n tu necesidad
.param Vcc = 5 ; Voltaje de referencia para la conversi�n
.param T = 1m  ; Periodo de la se�al de entrada y del reloj
*=============================================================================
* Calibration
*=============================================================================



*-----------------------------------------------------------------------------
*Libraries, Models and includes
*-----------------------------------------------------------------------------


*-----------------------------------------------------------------------------
*CIRCUIT
*-----------------------------------------------------------------------------
* Fuente de se�al anal�gica
;Vinput IN 0 SINE({FS/2} {FS/2} 1k)  ; Se�al senoidal con amplitud FS/2 y frecuencia de 1kHz
Vinput in 0 pwl(0 0 1m 0V 1.001m 2v 3m 2V  3.001m 0  5m 0V 6m 0v 6.001m 15v)

* Modelo de comportamiento del ADC de 4 bits
* Bit 3 (MSB) se activa si Vin >= FS * 8/16
B3 OUT[3] 0 V=if(V(in) >= {FS * 8 / 16}, 1, 0)

* Bit 2 se activa si Vin >= FS * 4/16, pero menos que el rango de bit 3
B2 OUT[2] 0 V=if(V(in) >= {FS * 4 / 16} & V(in) < {FS * 8 / 16}, 1, 0)

* Bit 1 se activa si Vin >= FS * 2/16, pero menos que el rango de bit 2 y 3
B1 OUT[1] 0 V=if(V(in) >= {FS * 2 / 16} & V(in) < {FS * 4 / 16}, 1, 0)

* Bit 0 (LSB) se activa si Vin >= FS * 1/16, pero menos que el rango de los bits superiores
B0 OUT[0] 0 V=if(V(in) >= {FS * 1 / 16} & V(in) < {FS * 2 / 16}, 1, 0)
* Resistores de carga en cada bit del bus;
R0 OUT[0] 0 1Meg
R1 OUT[1] 0 1Meg
R2 OUT[2] 0 1Meg
R3 OUT[3] 0 1Meg

* Fuente de reloj para la comparaci�n de bits
Vclk clk 0 PULSE(0 {Vcc} 0 1n 1n {T/2} {T})  ; Generador de reloj




;Vinput in 0 SINE(0 15 500) ;input
;Vinput in 0 pwl(0 0 1m 5V 4m 5V   6m 0V 7m 0v 7.001m 15v)
;Vinput in 0 pwl(1m 0 1.0001m 5v 2m 5v 2.001m 0v 3m 0v 3.001m 10v )

Vvdd Vdd 0 DC {p_Vfullscale}  ; Voltage full sacale

;if(x,y,z) If x > .5, then y else z


B0 out[0] 0 v={if(V(in)<{slope*1} ,0,if({V(in) <= {p_Vfullscale/((2*p_resolution)-1) * 1 & V(in)== {p_Vfullscale/((2*p_resolution)-1) } }
+| {V(in)=={p_Vfullscale/((2*p_resolution)-1) * 2}},1,0))}

;B1 out[1] 0 v={if(V(in)<{{V(in)>= {p_Vfullscale/((2*p_resolution)-1) * 2} }},0,if({V(in)>= {p_Vfullscale/((2*p_resolution)-1) * 3} } | {V(in)=={p_Vfullscale/((2*p_resolution)-1) * 4}},1,0))}



;Bout out 0 V =

*-----------------------------------------------------------------------------
*MEASUREMENTS
*-----------------------------------------------------------------------------


*-----------------------------------------------------------------------------
* SIMULATOR OPTIONS
*-----------------------------------------------------------------------------


*-----------------------------------------------------------------------------
* ANALYSIS
*-----------------------------------------------------------------------------
;.AC 	DEC 	10 	10 	10MEG
;.TRAN 	1US  	10m

.TRAN 10u 10m
.PROBE
.END
