*Half wave circuit with Diode
*------------------------------------------------------------------------------------------------------------------------------------------
*Circuit
*------------------------------------------------------------------------------------------------------------------------------------------
VS in	0	AC 1 SIN({p_offset} {p_ampl} {p_freq})
*------------------------------------------------------------------------------------------------------------------------------------------
D1 in	out	{Dmodel}
*D1 in	out	D
R1	out	0	{p_r1}
*------------------------------------------------------------------------------------------------------------------------------------------
*Models
*------------------------------------------------------------------------------------------------------------------------------------------
*.model D D
.model 1 ako:1N4148
.model 2 ako:1N5817
*------------------------------------------------------------------------------------------------------------------------------------------
*Standard library
*------------------------------------------------------------------------------------------------------------------------------------------
.lib C:\Users\jesse\AppData\Local\LTspice\lib\cmp\standard.dio
*------------------------------------------------------------------------------------------------------------------------------------------
*Parameters
*------------------------------------------------------------------------------------------------------------------------------------------
*.param p_r1	1k
.param p_r1		300; For 400mv, step 3
*Values of the wave
.param p_offset	0
.param p_ampl	1
.param p_freq	1k
*------------------------------------------------------------------------------------------------------------------------------------------
*mesures
*------------------------------------------------------------------------------------------------------------------------------------------
.meas	tran	Vout_max	MAX	V(out)
*------------------------------------------------------------------------------------------------------------------------------------------
* ANALYSIS
*------------------------------------------------------------------------------------------------------------------------------------------
.tran 10ms
.step param Dmodel list 1 2
*.step param p_r1 list 1k 5k
*Para calibracion de valores
*.step param p_r1  200 700 50 ;tener cuidado con la precision
.PLOT
.PROBE
.backanno;Annotate the Subcircuit Pin Names on Port Currents
.END
