adc_converter
*-----------------------------------------------------------------------------
*NOTES
*-----------------------------------------------------------------------------


*-----------------------------------------------------------------------------
*Parameters: User Input
*-----------------------------------------------------------------------------
.PARAM p_Vdd 15
.PARAM vthreshold 1

*=============================================================================
* Calibration
*=============================================================================



*-----------------------------------------------------------------------------
*Libraries, Models and includes
*-----------------------------------------------------------------------------
.LIB ADC_SAR.LIB

*-----------------------------------------------------------------------------
*CIRCUIT
*-----------------------------------------------------------------------------
Vin in 	0 PWL(0 0 20 20)
Vdd vdd 0 {p_Vdd}				; Fullscale

;.SUBCKT ADC_SAR_4bits in vdd vss out[3] out[2] out[1] out[0]
XDac_4bits in vdd 0 out1[3] out1[2] out1[1] out1[0] ADC_SAR_4bits

;.SUBCKT ADC_SAR_3bits in vdd vss out[3] out[2] out[1] out[0]
XDac_3bits in vdd 0 out2[2] out2[1] out2[0] ADC_SAR_3bits
*-----------------------------------------------------------------------------
*MEASUREMENTS
*-----------------------------------------------------------------------------
.INCLUDE ADC_SAR_MEASURMENTS.meas

*-----------------------------------------------------------------------------
* SIMULATOR OPTIONS
*-----------------------------------------------------------------------------


*-----------------------------------------------------------------------------
* ANALYSIS
*-----------------------------------------------------------------------------
;.AC 	DEC 	10 	10 	10MEG
;.TRAN 	1US  	10m
;.STEP PARAM p_Vdd list 5 15
.TRAN 10u 20
.PROBE
.END
