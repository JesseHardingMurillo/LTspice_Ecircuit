LowPassFilter
*-----------------------------------------------------------------------------
*NOTES
*-----------------------------------------------------------------------------
* This a LPF for replace with a step

*-----------------------------------------------------------------------------
*Libraries, Models and includes
*-----------------------------------------------------------------------------
.LIB LPF.LIB

*=============================================================================
* Calibration
*=============================================================================
.PARAM C 	5n
.PARAM fc 	5k


*-----------------------------------------------------------------------------
*CIRCUIT
*-----------------------------------------------------------------------------
*
VS	1	0	AC 1 SIN(0VOFF 1VPEAK 2KHZ)
*
;R1	1	2	{R}
;C1	2	0	{C}
XLPF 1 OUT LPF	PARAMS: C = {C}	fc = {fc}

*-----------------------------------------------------------------------------
* ANALYSIS
*-----------------------------------------------------------------------------
.AC 	DEC 	10 	10 	10MEG
;.TRAN 	1US  	10m
.PROBE
.END
